`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/04/2021 10:15:33 PM
// Design Name: 
// Module Name: PCsource_pkg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

package PCsource_pkg;

    localparam NEXT = 1'b0;
    localparam JUMP = 1'b1;
    
    // typedef enum logic { NEXT = 1'b0,
    //                      JUMP = 1'b1 } PCsource;
endpackage
